module pll_8_48(input clki, output clko);
	assign clko = clki;
endmodule
