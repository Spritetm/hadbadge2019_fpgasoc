module DP16KD (
    input ADA0,
    input ADA1,
    input ADA10,
    input ADA11,
    input ADA12,
    input ADA13,
    input ADA2,
    input ADA3,
    input ADA4,
    input ADA5,
    input ADA6,
    input ADA7,
    input ADA8,
    input ADA9,
    input ADB0,
    input ADB1,
    input ADB10,
    input ADB11,
    input ADB12,
    input ADB13,
    input ADB2,
    input ADB3,
    input ADB4,
    input ADB5,
    input ADB6,
    input ADB7,
    input ADB8,
    input ADB9,
    input CEA,
    input CEB,
    input CLKA,
    input CLKB,
    input DIA0,
    input DIA1,
    input DIA10,
    input DIA11,
    input DIA12,
    input DIA13,
    input DIA14,
    input DIA15,
    input DIA16,
    input DIA17,
    input DIA2,
    input DIA3,
    input DIA4,
    input DIA5,
    input DIA6,
    input DIA7,
    input DIA8,
    input DIA9,
    input DIB0,
    input DIB1,
    input DIB10,
    input DIB11,
    input DIB12,
    input DIB13,
    input DIB14,
    input DIB15,
    input DIB16,
    input DIB17,
    input DIB2,
    input DIB3,
    input DIB4,
    input DIB5,
    input DIB6,
    input DIB7,
    input DIB8,
    input DIB9,
    output DOA0,
    output DOA1,
    output DOA10,
    output DOA11,
    output DOA12,
    output DOA13,
    output DOA14,
    output DOA15,
    output DOA16,
    output DOA17,
    output DOA2,
    output DOA3,
    output DOA4,
    output DOA5,
    output DOA6,
    output DOA7,
    output DOA8,
    output DOA9,
    output DOB0,
    output DOB1,
    output DOB10,
    output DOB11,
    output DOB12,
    output DOB13,
    output DOB14,
    output DOB15,
    output DOB16,
    output DOB17,
    output DOB2,
    output DOB3,
    output DOB4,
    output DOB5,
    output DOB6,
    output DOB7,
    output DOB8,
    output DOB9,
    input OCEA,
    input OCEB,
    input RSTA,
    input RSTB,
    input WEA,
    input WEB
  );

    parameter CLKAMUX = "CLKA";
    parameter CLKBMUX = "CLKB";
    parameter DATA_WIDTH_A = 32'd4;
    parameter DATA_WIDTH_B = 32'd4;
    parameter GSR = "DISABLED";
    parameter INITVAL_00 = 320'h13020092980c29619aa305a2202e0b0b0df104560dee61fcad096d212cb7060360d8e61e89e15698;
    parameter INITVAL_01 = 320'h008e50646a0fe9d0c0b5106f60f8b4072e501cf6178e6174b3162b515cbc1846a104ff01cd106e31;
    parameter INITVAL_02 = 320'h0e6fa172fb1c4ae096280a8210b65c03ec71b6bf08a3c01470156851fea5028fc1a4330888f0ce52;
    parameter INITVAL_03 = 320'h100f00d837106720b8d20d04d1b4be1a4ab16e9504a2113a421d8831a4290e84717c1b0fe0418e3f;
    parameter INITVAL_04 = 320'h0e03d020971509103409176d81a6e0006960ee360904909c0e00ceb13a5405e851227206276062cf;
    parameter INITVAL_05 = 320'h116801d4a503c600b2e80f4740548f1281912a0a1e477034610ceee1280b128d5084bf1707502413;
    parameter INITVAL_06 = 320'h16aeb09ea2112bb098a8036a714a1202cdc1609b0f85813c08114130b06d0bc391f0a219e7f1ca6f;
    parameter INITVAL_07 = 320'h00e1f1467113c8c040aa044721908a148071f2d01cad60c0811fa140ea10194060224900ed10a6fa;
    parameter INITVAL_08 = 320'h0e4c61a02f0c0320a82d0c437024670424a0b4e8070ae076fd04a190fca71800b1249d1f43f02c09;
    parameter INITVAL_09 = 320'h1e08003a42176a21e6cc1241f1a239048090764e0f80d0983b1d07c054af038bb1a0de0789207efb;
    parameter INITVAL_0A = 320'h19c4b120451988618e2806ea703ed00b2d11ca1801604106fa14e51168c7176470f20011816062a1;
    parameter INITVAL_0B = 320'h04837066fa0543c00263100a40a44209a4b166b50da9601405006ff16cac1127717e0a0167f14c3b;
    parameter INITVAL_0C = 320'h19ee607cc60f0ec1564406c9118e52172410e89303cf4150e8058e10f4e51a42518e9108a611b612;
    parameter INITVAL_0D = 320'h0b0790d826168a30f0540766501e210a213006bd1fcdd026f51f2951d66507c63084d30c8ce06856;
    parameter INITVAL_0E = 320'h0dacf1d4a7110cc09ed30ac8c1c2370c48102aba0b8c41fe820066f0b42f16a021f6fb12eb50003d;
    parameter INITVAL_0F = 320'h18cd215e2f1047e0284702e38128890207b0ee140fc760a08c1880a0e8f70c8ed1d46d17a711f055;
    parameter INITVAL_10 = 320'h1e89e1a671046c50803f008fc0d09d018df1d0de196aa098cd1162b0a029012611321019c4616a93;
    parameter INITVAL_11 = 320'h1e4ab18edf112251ee4908e510a62007016146b60466b05a491d610032041a8731ea2e0a2b61c0b0;
    parameter INITVAL_12 = 320'h0aea2098b21decc130230842d19a180742f0967b098c116eb419e381382b1c85405c90094511044a;
    parameter INITVAL_13 = 320'h0b2100d06c10e75122020028c06c710709a1e2181aea60522a0181208a86078e40a6790e21d04a35;
    parameter INITVAL_14 = 320'h150011943313c021b80a16cee1205c092950969c16e5f0ca201e0851ecf41faef1789e00aae0ee35;
    parameter INITVAL_15 = 320'h1882d19c551c4c91e43514c380b04219c2803cb016aa81b61818c1405a8213a440523a0f0ce0f400;
    parameter INITVAL_16 = 320'h092721ca2d15038000f8168570f4551fc08056121c86a156670843713c0f08c560b0201b8e30cc2d;
    parameter INITVAL_17 = 320'h10e0d0d075148de05c6813af30c6e0182ec102e00642707c971b4da04a5f00af0026b90408b1944b;
    parameter INITVAL_18 = 320'h16ca206eb41e4960aa691501d006de0d2890e6ff16c4c0549a1dc380ae9d0ac4d186630842b0d0cc;
    parameter INITVAL_19 = 320'h0727a0fabc10cfc1c618124421c29d0b882112d90c41618018194d8086ac146221a0b704af50ce95;
    parameter INITVAL_1A = 320'h1068213253190991b2d91c05107ecf11c890e03014ecd156321c4921924c132581d69a196fe01287;
    parameter INITVAL_1B = 320'h18e4c19af409a5c116f71f49c1786c17e0009c080e64d086a30ea241cceb0d69119a581b0ea19610;
    parameter INITVAL_1C = 320'h19e6503835088c409e4713eba126c213ac61ea6a038f41401800e911fafb0be4f1280313ccf12438;
    parameter INITVAL_1D = 320'h02c031961a0f60101e75024c013e6f166971e4601d0df1e01a160b116e3c0acb5064b6166b3168a9;
    parameter INITVAL_1E = 320'h1b02d1b2a712a9718afa170a81863013ce61a006098f01e48f0b26a01c1d1407c190e703e7c18870;
    parameter INITVAL_1F = 320'h15c2d1aa661cc421247517ad517c3c134270848c056481bc740504005c41158ca0fc980b02f1501e;
    parameter INITVAL_20 = 320'h0f4bf1a283076d81f8fa0163310875006c61e8091d035186b80060800c3918ec010205116b61083f;
    parameter INITVAL_21 = 320'h09ac308cb5152391b4490f8970cced18a9f0d4991240d0a69700a781ac1d158830f80c038f618cba;
    parameter INITVAL_22 = 320'h166aa08e0e1d8ca0821a0862815c5f0068a07c8715af608a271f0bc1543e1f4560d2ae1e4671a480;
    parameter INITVAL_23 = 320'h188241022503214168450b277140e5094fd1b05d0dee011ede130161ea4d190ae1c8d00e07816e93;
    parameter INITVAL_24 = 320'h0b28e14cb902e951049f152fc196bf050f708618174f0108070ac20018b708c3b19e8b0d6951d2a7;
    parameter INITVAL_25 = 320'h15811036f20529013ee319eaf0567a0b6171cc5e13a2506a321dab80c8ee1ae0c150c711e7a0169f;
    parameter INITVAL_26 = 320'h0246f0dc891d8871e0760ca4c088271e0851ca2b0881b0149f114591d46412a54048bc1ea320cccf;
    parameter INITVAL_27 = 320'h19a5200e39174441807805a6e1f2cd17abd012bc092750a4c100602152cd0e4e90da3108c81148a8;
    parameter INITVAL_28 = 320'h170a01ee6319e6114a6914aa2110d0196780fcb2156961201512c930de4100a41176250c4b800cea;
    parameter INITVAL_29 = 320'h1a87910cbc0aa17042e101a2d134e21969116e8801afb1684e0beb4062c913063110f9086ef070f6;
    parameter INITVAL_2A = 320'h1b4be1ee62106dd1269118eda11c3c0d49b0782f1aefe086f001ad9028f01d2fd08a281d6251b401;
    parameter INITVAL_2B = 320'h00a331aa2618e53106bf0021f1bcb204ce10d8680f8d50b4c10801615c8a150dd0e4f31f6dc1004d;
    parameter INITVAL_2C = 320'h164c4074831263c112d411e2b04c141beb80a6bb016fd0225c0d6b9082961749a1aacb1bc451de5f;
    parameter INITVAL_2D = 320'h1eeda012831ecd80da92034ca0348d0ce770664d14ac512a6f0c4c2116c705e4c00e94086710be28;
    parameter INITVAL_2E = 320'h00a1405cde0d67b0fa7d0cc031b8931ae841a60c0ce8d0462e076851ec121a6d90768a0aa4d18eb0;
    parameter INITVAL_2F = 320'h0ca4e1b2630a650124a8048be04e601d83204c730862901c57166e71b45a0c0e2144821ecd21363d;
    parameter INITVAL_30 = 320'h132f9008c3176d81de24046461ead00a8ca01c750062c064fe1fe5a0ce2f1d2f70429a1f20319077;
    parameter INITVAL_31 = 320'h1ce23076bf0b2e30bc2b0ccbb0e8f9054150ce691f674196201001a02a520d4f4000fe16089014c6;
    parameter INITVAL_32 = 320'h0d864040a606cab1beba0fe680f65d0464b134e21b6351c06d0a0a11682e0e85e00e6d08e9f074f0;
    parameter INITVAL_33 = 320'h1c06012ede04e7a0a637056be01807144fb076b31d06a180160caa702ce1018421c2f10846c1521c;
    parameter INITVAL_34 = 320'h124b0092a50da20110d107cec040c912a0717a3e02c1b166de1c2f6094ca0cc6e14efa0da9e19e54;
    parameter INITVAL_35 = 320'h1a2d91f89e14c3c0e6640bc011c074198a10700f1084a040180087905813166a91ba8b018f4056e5;
    parameter INITVAL_36 = 320'h0beb60ca390de8f03aff0a21a0fa30072fe12e6f078901ccc11f8a903c8208e51010df0426c09a53;
    parameter INITVAL_37 = 320'h122540c4fd1481e05235040511743e10afd1b07f05eee024cc16a681ea3d1c4f80c0461cce40c094;
    parameter INITVAL_38 = 320'h0c8d81ecd0056b60445909cf41dab91249207ad4064951d2aa104a5068d9136a3038a603e561beef;
    parameter INITVAL_39 = 320'h05a18128e61742a060d906e240aa4f086a81484a19aaf16af01c62e06abe0e6920123e1c44b1c88a;
    parameter INITVAL_3A = 320'h0ec4c018a217a6e0f0e815e2c1ce74192521bc49178651e6f31162e086b414c7c0829406e2418e4f;
    parameter INITVAL_3B = 320'h016461b8a40c40b086a50a2100c8a708a9808a050722a0122d13a9c19e821f6f70d6490683e1dab6;
    parameter INITVAL_3C = 320'h1769e0f2611bc951889d0eadd12eb60b6990222b166771069a0fc6c0d89d01ec2198ce0b0d402224;
    parameter INITVAL_3D = 320'h01ade07c950c8f81fc5413a2d0d81a1d4561c6ac086a716e530f2f113e4d1425f142111440e128ac;
    parameter INITVAL_3E = 320'h1004d072091de16056b81208b1a09a0d07910a61150fd046720d08d17ea5062c51c43018a8f04489;
    parameter INITVAL_3F = 320'h0103918ab0108961ced31ea841f8f60803907c251c6a70cc26170e716a5d1aec00387f18692060e3;
    parameter WRITEMODE_A = "READBEFOREWRITE";
    parameter WRITEMODE_B = "READBEFOREWRITE";


	wire [13:0] ADA;
	assign ADA = {ADA13, ADA12, ADA11, ADA10, ADA9, ADA8, ADA7, ADA6, ADA5, ADA4, ADA3, ADA2, ADA1, ADA0};
	wire [13:0] ADB;
	assign ADB = {ADB13, ADB12, ADB11, ADB10, ADB9, ADB8, ADB7, ADB6, ADB5, ADB4, ADB3, ADB2, ADB1, ADB0};
	wire [17:0] DIA;
	assign DIA = {DIA17, DIA16, DIA15, DIA14, DIA13, DIA12, DIA11, DIA10, DIA9, DIA8, DIA7, DIA6, DIA5, DIA4, DIA3, DIA2, DIA1, DIA0};
	wire [17:0] DIB;
	assign DIB = {DIB17, DIB16, DIB15, DIB14, DIB13, DIB12, DIB11, DIB10, DIB9, DIB8, DIB7, DIB6, DIB5, DIB4, DIB3, DIB2, DIB1, DIB0};
	wire [17:0] DOA;
	assign {DOA17, DOA16, DOA15, DOA14, DOA13, DOA12, DOA11, DOA10, DOA9, DOA8, DOA7, DOA6, DOA5, DOA4, DOA3, DOA2, DOA1, DOA0}=DOA;
	wire [17:0] DOB;
	assign {DOB17, DOB16, DOB15, DOB14, DOB13, DOB12, DOB11, DOB10, DOB9, DOB8, DOB7, DOB6, DOB5, DOB4, DOB3, DOB2, DOB1, DOB0}=DOB;


endmodule