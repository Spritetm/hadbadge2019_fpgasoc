

module vid_tilemapmem (DataInA, DataInB, AddressA, AddressB, ClockA, 
    ClockB, ClockEnA, ClockEnB, WrA, WrB, ResetA, ResetB, QA, QB);
    input wire [17:0] DataInA;
    input wire [17:0] DataInB;
    input wire [11:0] AddressA;
    input wire [11:0] AddressB;
    input wire ClockA;
    input wire ClockB;
    input wire ClockEnA;
    input wire ClockEnB;
    input wire WrA;
    input wire WrB;
    input wire ResetA;
    input wire ResetB;
    output wire [17:0] QA;
    output wire [17:0] QB;

wire [17:0] qa1;
wire [17:0] qb1;
wire [17:0] qa2;
wire [17:0] qb2;

vid_tilemapmem_2kx18_ecp5 mem1(
	.DataInA(DataInA),
	.DataInB(DataInB),
	.AddressA(AddressA[10:0]),
	.AddressB(AddressB[10:0]),
	.ClockA(ClockA),
	.ClockB(ClockB),
	.ClockEnA(ClockEnA),
	.ClockEnB(ClockEnB),
	.WrA(WrA & (~AddressA[11])),
	.WrB(WrB & (~AddressB[11])),
	.ResetA(ResetA),
	.ResetB(ResetB),
	.QA(qa1),
	.QB(qb1)
);

vid_tilemapmem_2kx18_ecp5 mem2(
	.DataInA(DataInA),
	.DataInB(DataInB),
	.AddressA(AddressA[10:0]),
	.AddressB(AddressB[10:0]),
	.ClockA(ClockA),
	.ClockB(ClockB),
	.ClockEnA(ClockEnA),
	.ClockEnB(ClockEnB),
	.WrA(WrA & AddressA[11]),
	.WrB(WrB & AddressB[11]),
	.ResetA(ResetA),
	.ResetB(ResetB),
	.QA(qa2),
	.QB(qb2)
);

reg addra_reg;
always @(posedge ClockA) begin
	addra_reg <= AddressA[11];
end
reg addrb_reg;
always @(posedge ClockB) begin
	addrb_reg <= AddressB[11];
end

assign QA = addra_reg ? qa2 : qa1;
assign QB = addrb_reg ? qb2 : qb1;

endmodule


/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.10.2.115.2 */
/* Module Version: 7.5 */
/* /home/jeroen/diamond/ispfpga/bin/lin64/scuba -w -n vid_tilemem_2kx18 -lang verilog -synth lse -bus_exp 7 -bb -arch sa5p00 -type bram -wp 11 -rp 1010 -data_width 18 -rdata_width 18 -num_rows 2048 -outdataA REGISTERED -outdataB REGISTERED -cascade -1 -resetmode SYNC -sync_reset -mem_init0 -writemodeA NORMAL -writemodeB NORMAL -fdc /tmp/test/vid_tilemem/vid_tilemem_2kx18/vid_tilemem_2kx18.fdc  */
/* Sun Sep 29 22:16:40 2019 */

`timescale 1 ns / 1 ps
module vid_tilemapmem_2kx18_ecp5 (DataInA, DataInB, AddressA, AddressB, ClockA, 
    ClockB, ClockEnA, ClockEnB, WrA, WrB, ResetA, ResetB, QA, QB)/* synthesis NGD_DRC_MASK=1 */;
    input wire [17:0] DataInA;
    input wire [17:0] DataInB;
    input wire [10:0] AddressA;
    input wire [10:0] AddressB;
    input wire ClockA;
    input wire ClockB;
    input wire ClockEnA;
    input wire ClockEnB;
    input wire WrA;
    input wire WrB;
    input wire ResetA;
    input wire ResetB;
    output wire [17:0] QA;
    output wire [17:0] QB;

    wire scuba_vhi;
    wire scuba_vlo;
    assign scuba_vhi = 1;
    assign scuba_vlo = 0;

//    defparam vid_tilemem_2kx18_0_0_1.INIT_DATA = "STATIC" ;
    defparam vid_tilemem_2kx18_0_0_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_0_1.CSDECODE_B = "0b000" ;
    defparam vid_tilemem_2kx18_0_0_1.CSDECODE_A = "0b000" ;
    defparam vid_tilemem_2kx18_0_0_1.WRITEMODE_B = "NORMAL" ;
    defparam vid_tilemem_2kx18_0_0_1.WRITEMODE_A = "NORMAL" ;
    defparam vid_tilemem_2kx18_0_0_1.GSR = "ENABLED" ;
    defparam vid_tilemem_2kx18_0_0_1.RESETMODE = "SYNC" ;
    defparam vid_tilemem_2kx18_0_0_1.REGMODE_B = "OUTREG" ;
    defparam vid_tilemem_2kx18_0_0_1.REGMODE_A = "OUTREG" ;
    defparam vid_tilemem_2kx18_0_0_1.DATA_WIDTH_B = 9 ;
    defparam vid_tilemem_2kx18_0_0_1.DATA_WIDTH_A = 9 ;
    DP16KD vid_tilemem_2kx18_0_0_1 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(DataInA[8]), 
        .DIA7(DataInA[7]), .DIA6(DataInA[6]), .DIA5(DataInA[5]), .DIA4(DataInA[4]), 
        .DIA3(DataInA[3]), .DIA2(DataInA[2]), .DIA1(DataInA[1]), .DIA0(DataInA[0]), 
        .ADA13(AddressA[10]), .ADA12(AddressA[9]), .ADA11(AddressA[8]), 
        .ADA10(AddressA[7]), .ADA9(AddressA[6]), .ADA8(AddressA[5]), .ADA7(AddressA[4]), 
        .ADA6(AddressA[3]), .ADA5(AddressA[2]), .ADA4(AddressA[1]), .ADA3(AddressA[0]), 
        .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(DataInB[8]), 
        .DIB7(DataInB[7]), .DIB6(DataInB[6]), .DIB5(DataInB[5]), .DIB4(DataInB[4]), 
        .DIB3(DataInB[3]), .DIB2(DataInB[2]), .DIB1(DataInB[1]), .DIB0(DataInB[0]), 
        .ADB13(AddressB[10]), .ADB12(AddressB[9]), .ADB11(AddressB[8]), 
        .ADB10(AddressB[7]), .ADB9(AddressB[6]), .ADB8(AddressB[5]), .ADB7(AddressB[4]), 
        .ADB6(AddressB[3]), .ADB5(AddressB[2]), .ADB4(AddressB[1]), .ADB3(AddressB[0]), 
        .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(QA[8]), .DOA7(QA[7]), 
        .DOA6(QA[6]), .DOA5(QA[5]), .DOA4(QA[4]), .DOA3(QA[3]), .DOA2(QA[2]), 
        .DOA1(QA[1]), .DOA0(QA[0]), .DOB17(), .DOB16(), .DOB15(), .DOB14(), 
        .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), .DOB8(QB[8]), .DOB7(QB[7]), 
        .DOB6(QB[6]), .DOB5(QB[5]), .DOB4(QB[4]), .DOB3(QB[3]), .DOB2(QB[2]), 
        .DOB1(QB[1]), .DOB0(QB[0]))
             /* synthesis MEM_LPC_FILE="vid_tilemem_2kx18.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;


//    defparam vid_tilemem_2kx18_0_1_0.INIT_DATA = "STATIC" ;
    defparam vid_tilemem_2kx18_0_1_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam vid_tilemem_2kx18_0_1_0.CSDECODE_B = "0b000" ;
    defparam vid_tilemem_2kx18_0_1_0.CSDECODE_A = "0b000" ;
    defparam vid_tilemem_2kx18_0_1_0.WRITEMODE_B = "NORMAL" ;
    defparam vid_tilemem_2kx18_0_1_0.WRITEMODE_A = "NORMAL" ;
    defparam vid_tilemem_2kx18_0_1_0.GSR = "ENABLED" ;
    defparam vid_tilemem_2kx18_0_1_0.RESETMODE = "SYNC" ;
    defparam vid_tilemem_2kx18_0_1_0.REGMODE_B = "OUTREG" ;
    defparam vid_tilemem_2kx18_0_1_0.REGMODE_A = "OUTREG" ;
    defparam vid_tilemem_2kx18_0_1_0.DATA_WIDTH_B = 9 ;
    defparam vid_tilemem_2kx18_0_1_0.DATA_WIDTH_A = 9 ;
    DP16KD vid_tilemem_2kx18_0_1_0 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(DataInA[17]), 
        .DIA7(DataInA[16]), .DIA6(DataInA[15]), .DIA5(DataInA[14]), .DIA4(DataInA[13]), 
        .DIA3(DataInA[12]), .DIA2(DataInA[11]), .DIA1(DataInA[10]), .DIA0(DataInA[9]), 
        .ADA13(AddressA[10]), .ADA12(AddressA[9]), .ADA11(AddressA[8]), 
        .ADA10(AddressA[7]), .ADA9(AddressA[6]), .ADA8(AddressA[5]), .ADA7(AddressA[4]), 
        .ADA6(AddressA[3]), .ADA5(AddressA[2]), .ADA4(AddressA[1]), .ADA3(AddressA[0]), 
        .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(DataInB[17]), 
        .DIB7(DataInB[16]), .DIB6(DataInB[15]), .DIB5(DataInB[14]), .DIB4(DataInB[13]), 
        .DIB3(DataInB[12]), .DIB2(DataInB[11]), .DIB1(DataInB[10]), .DIB0(DataInB[9]), 
        .ADB13(AddressB[10]), .ADB12(AddressB[9]), .ADB11(AddressB[8]), 
        .ADB10(AddressB[7]), .ADB9(AddressB[6]), .ADB8(AddressB[5]), .ADB7(AddressB[4]), 
        .ADB6(AddressB[3]), .ADB5(AddressB[2]), .ADB4(AddressB[1]), .ADB3(AddressB[0]), 
        .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(QA[17]), 
        .DOA7(QA[16]), .DOA6(QA[15]), .DOA5(QA[14]), .DOA4(QA[13]), .DOA3(QA[12]), 
        .DOA2(QA[11]), .DOA1(QA[10]), .DOA0(QA[9]), .DOB17(), .DOB16(), 
        .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), .DOB10(), .DOB9(), 
        .DOB8(QB[17]), .DOB7(QB[16]), .DOB6(QB[15]), .DOB5(QB[14]), .DOB4(QB[13]), 
        .DOB3(QB[12]), .DOB2(QB[11]), .DOB1(QB[10]), .DOB0(QB[9]))
             /* synthesis MEM_LPC_FILE="vid_tilemem_2kx18.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;



    // exemplar begin
    // exemplar attribute vid_tilemem_2kx18_0_0_1 MEM_LPC_FILE vid_tilemem_2kx18.lpc
    // exemplar attribute vid_tilemem_2kx18_0_0_1 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute vid_tilemem_2kx18_0_1_0 MEM_LPC_FILE vid_tilemem_2kx18.lpc
    // exemplar attribute vid_tilemem_2kx18_0_1_0 MEM_INIT_FILE INIT_ALL_0s
    // exemplar end

endmodule
