
`timescale 1 ns / 1 ps
module vid_tilemem (DataInA, DataInB, AddressA, AddressB, ClockA, 
    ClockB, ClockEnA, ClockEnB, WrA, WrB, ResetA, ResetB, QA, QB)/* synthesis NGD_DRC_MASK=1 */;
    input wire [31:0] DataInA;
    input wire [31:0] DataInB;
    input wire [13:0] AddressA;
    input wire [13:0] AddressB;
    input wire ClockA;
    input wire ClockB;
    input wire ClockEnA;
    input wire ClockEnB;
    input wire WrA;
    input wire WrB;
    input wire ResetA;
    input wire ResetB;
    output wire [31:0] QA;
    output wire [31:0] QB;

    wire scuba_vhi;
    wire scuba_vlo;

    //VHI scuba_vhi_inst (.Z(scuba_vhi));
	assign scuba_vhi = 1;
	assign scuba_vlo = 0;

//    defparam tilemem_ecp5_inst_0_0_31.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_0_31.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_0_31.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_0_31.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_0_31.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_0_31.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_0_31.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_0_31.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_0_31.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_0_31.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_0_31.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_0_31.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_0_31 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[0]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[0]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[0]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[0]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_1_30.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_1_30.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_1_30.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_1_30.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_1_30.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_1_30.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_1_30.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_1_30.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_1_30.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_1_30.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_1_30.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_1_30.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_1_30 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[1]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[1]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[1]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[1]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_2_29.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_2_29.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_2_29.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_2_29.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_2_29.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_2_29.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_2_29.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_2_29.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_2_29.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_2_29.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_2_29.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_2_29.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_2_29 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[2]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[2]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[2]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[2]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_3_28.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_3_28.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_3_28.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_3_28.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_3_28.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_3_28.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_3_28.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_3_28.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_3_28.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_3_28.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_3_28.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_3_28.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_3_28 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[3]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[3]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[3]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[3]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_4_27.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_4_27.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_4_27.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_4_27.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_4_27.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_4_27.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_4_27.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_4_27.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_4_27.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_4_27.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_4_27.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_4_27.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_4_27 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[4]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[4]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[4]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[4]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_5_26.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_5_26.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_5_26.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_5_26.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_5_26.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_5_26.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_5_26.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_5_26.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_5_26.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_5_26.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_5_26.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_5_26.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_5_26 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[5]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[5]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[5]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[5]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_6_25.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_6_25.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_6_25.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_6_25.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_6_25.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_6_25.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_6_25.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_6_25.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_6_25.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_6_25.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_6_25.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_6_25.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_6_25 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[6]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[6]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[6]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[6]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_7_24.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_7_24.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_7_24.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_7_24.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_7_24.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_7_24.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_7_24.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_7_24.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_7_24.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_7_24.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_7_24.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_7_24.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_7_24 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[7]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[7]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[7]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[7]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_8_23.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_8_23.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_8_23.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_8_23.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_8_23.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_8_23.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_8_23.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_8_23.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_8_23.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_8_23.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_8_23.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_8_23.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_8_23 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[8]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[8]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[8]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[8]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_9_22.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_9_22.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_9_22.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_9_22.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_9_22.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_9_22.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_9_22.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_9_22.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_9_22.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_9_22.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_9_22.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_9_22.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_9_22 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[9]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[9]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[9]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[9]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_10_21.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_10_21.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_10_21.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_10_21.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_10_21.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_10_21.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_10_21.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_10_21.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_10_21.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_10_21.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_10_21.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_10_21.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_10_21 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[10]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[10]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[10]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[10]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_11_20.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_11_20.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_11_20.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_11_20.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_11_20.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_11_20.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_11_20.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_11_20.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_11_20.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_11_20.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_11_20.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_11_20.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_11_20 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[11]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[11]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[11]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[11]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_12_19.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_12_19.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_12_19.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_12_19.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_12_19.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_12_19.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_12_19.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_12_19.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_12_19.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_12_19.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_12_19.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_12_19.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_12_19 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[12]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[12]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[12]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[12]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_13_18.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_13_18.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_13_18.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_13_18.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_13_18.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_13_18.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_13_18.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_13_18.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_13_18.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_13_18.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_13_18.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_13_18.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_13_18 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[13]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[13]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[13]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[13]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_14_17.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_14_17.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_14_17.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_14_17.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_14_17.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_14_17.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_14_17.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_14_17.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_14_17.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_14_17.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_14_17.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_14_17.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_14_17 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[14]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[14]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[14]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[14]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_15_16.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_15_16.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_15_16.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_15_16.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_15_16.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_15_16.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_15_16.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_15_16.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_15_16.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_15_16.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_15_16.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_15_16.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_15_16 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[15]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[15]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[15]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[15]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_16_15.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_16_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_16_15.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_16_15.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_16_15.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_16_15.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_16_15.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_16_15.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_16_15.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_16_15.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_16_15.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_16_15.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_16_15 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[16]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[16]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[16]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[16]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_17_14.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_17_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_17_14.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_17_14.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_17_14.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_17_14.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_17_14.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_17_14.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_17_14.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_17_14.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_17_14.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_17_14.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_17_14 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[17]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[17]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[17]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[17]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_18_13.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_18_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_18_13.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_18_13.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_18_13.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_18_13.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_18_13.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_18_13.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_18_13.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_18_13.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_18_13.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_18_13.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_18_13 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[18]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[18]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[18]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[18]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_19_12.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_19_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_19_12.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_19_12.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_19_12.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_19_12.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_19_12.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_19_12.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_19_12.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_19_12.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_19_12.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_19_12.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_19_12 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[19]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[19]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[19]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[19]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_20_11.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_20_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_20_11.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_20_11.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_20_11.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_20_11.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_20_11.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_20_11.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_20_11.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_20_11.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_20_11.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_20_11.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_20_11 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[20]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[20]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[20]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[20]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_21_10.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_21_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_21_10.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_21_10.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_21_10.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_21_10.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_21_10.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_21_10.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_21_10.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_21_10.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_21_10.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_21_10.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_21_10 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[21]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[21]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[21]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[21]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_22_9.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_22_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_22_9.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_22_9.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_22_9.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_22_9.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_22_9.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_22_9.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_22_9.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_22_9.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_22_9.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_22_9.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_22_9 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[22]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[22]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[22]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[22]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_23_8.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_23_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_23_8.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_23_8.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_23_8.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_23_8.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_23_8.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_23_8.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_23_8.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_23_8.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_23_8.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_23_8.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_23_8 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[23]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[23]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[23]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[23]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_24_7.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_24_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_24_7.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_24_7.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_24_7.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_24_7.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_24_7.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_24_7.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_24_7.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_24_7.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_24_7.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_24_7.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_24_7 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[24]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[24]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[24]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[24]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_25_6.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_25_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_25_6.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_25_6.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_25_6.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_25_6.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_25_6.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_25_6.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_25_6.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_25_6.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_25_6.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_25_6.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_25_6 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[25]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[25]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[25]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[25]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_26_5.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_26_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_26_5.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_26_5.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_26_5.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_26_5.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_26_5.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_26_5.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_26_5.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_26_5.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_26_5.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_26_5.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_26_5 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[26]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[26]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[26]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[26]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_27_4.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_27_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_27_4.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_27_4.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_27_4.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_27_4.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_27_4.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_27_4.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_27_4.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_27_4.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_27_4.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_27_4.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_27_4 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[27]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[27]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[27]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[27]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_28_3.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_28_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_28_3.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_28_3.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_28_3.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_28_3.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_28_3.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_28_3.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_28_3.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_28_3.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_28_3.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_28_3.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_28_3 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[28]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[28]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[28]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[28]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_29_2.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_29_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_29_2.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_29_2.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_29_2.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_29_2.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_29_2.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_29_2.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_29_2.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_29_2.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_29_2.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_29_2.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_29_2 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[29]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[29]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[29]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[29]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

//    defparam tilemem_ecp5_inst_0_30_1.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_30_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_30_1.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_30_1.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_30_1.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_30_1.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_30_1.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_30_1.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_30_1.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_30_1.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_30_1.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_30_1.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_30_1 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[30]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[30]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[30]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[30]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;

    //VLO scuba_vlo_inst (.Z(scuba_vlo));

//    defparam tilemem_ecp5_inst_0_31_0.INIT_DATA = "STATIC" ;
    defparam tilemem_ecp5_inst_0_31_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_3F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_38 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_37 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_36 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_35 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_34 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_33 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_32 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_31 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_30 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_2F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_2E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_2D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_2C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_2B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_2A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_29 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_28 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_27 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_26 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_25 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_24 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_23 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_22 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_21 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_20 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam tilemem_ecp5_inst_0_31_0.CSDECODE_B = "0b000" ;
    defparam tilemem_ecp5_inst_0_31_0.CSDECODE_A = "0b000" ;
    defparam tilemem_ecp5_inst_0_31_0.WRITEMODE_B = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_31_0.WRITEMODE_A = "NORMAL" ;
    defparam tilemem_ecp5_inst_0_31_0.GSR = "ENABLED" ;
    defparam tilemem_ecp5_inst_0_31_0.RESETMODE = "SYNC" ;
    defparam tilemem_ecp5_inst_0_31_0.REGMODE_B = "NOREG" ;
    defparam tilemem_ecp5_inst_0_31_0.REGMODE_A = "NOREG" ;
    defparam tilemem_ecp5_inst_0_31_0.DATA_WIDTH_B = 1 ;
    defparam tilemem_ecp5_inst_0_31_0.DATA_WIDTH_A = 1 ;
    DP16KD tilemem_ecp5_inst_0_31_0 (.DIA17(scuba_vlo), .DIA16(scuba_vlo), 
        .DIA15(scuba_vlo), .DIA14(scuba_vlo), .DIA13(scuba_vlo), .DIA12(scuba_vlo), 
        .DIA11(scuba_vlo), .DIA10(scuba_vlo), .DIA9(scuba_vlo), .DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(DataInA[31]), 
        .ADA13(AddressA[13]), .ADA12(AddressA[12]), .ADA11(AddressA[11]), 
        .ADA10(AddressA[10]), .ADA9(AddressA[9]), .ADA8(AddressA[8]), .ADA7(AddressA[7]), 
        .ADA6(AddressA[6]), .ADA5(AddressA[5]), .ADA4(AddressA[4]), .ADA3(AddressA[3]), 
        .ADA2(AddressA[2]), .ADA1(AddressA[1]), .ADA0(AddressA[0]), .CEA(ClockEnA), 
        .OCEA(ClockEnA), .CLKA(ClockA), .WEA(WrA), .CSA2(scuba_vlo), .CSA1(scuba_vlo), 
        .CSA0(scuba_vlo), .RSTA(ResetA), .DIB17(scuba_vlo), .DIB16(scuba_vlo), 
        .DIB15(scuba_vlo), .DIB14(scuba_vlo), .DIB13(scuba_vlo), .DIB12(scuba_vlo), 
        .DIB11(scuba_vlo), .DIB10(scuba_vlo), .DIB9(scuba_vlo), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(DataInB[31]), 
        .ADB13(AddressB[13]), .ADB12(AddressB[12]), .ADB11(AddressB[11]), 
        .ADB10(AddressB[10]), .ADB9(AddressB[9]), .ADB8(AddressB[8]), .ADB7(AddressB[7]), 
        .ADB6(AddressB[6]), .ADB5(AddressB[5]), .ADB4(AddressB[4]), .ADB3(AddressB[3]), 
        .ADB2(AddressB[2]), .ADB1(AddressB[1]), .ADB0(AddressB[0]), .CEB(ClockEnB), 
        .OCEB(ClockEnB), .CLKB(ClockB), .WEB(WrB), .CSB2(scuba_vlo), .CSB1(scuba_vlo), 
        .CSB0(scuba_vlo), .RSTB(ResetB), .DOA17(), .DOA16(), .DOA15(), .DOA14(), 
        .DOA13(), .DOA12(), .DOA11(), .DOA10(), .DOA9(), .DOA8(), .DOA7(), 
        .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(QA[31]), 
        .DOB17(), .DOB16(), .DOB15(), .DOB14(), .DOB13(), .DOB12(), .DOB11(), 
        .DOB10(), .DOB9(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(QB[31]))
             /* synthesis MEM_LPC_FILE="tilemem_ecp5_inst.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;



    // exemplar begin
    // exemplar attribute tilemem_ecp5_inst_0_0_31 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_0_31 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_1_30 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_1_30 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_2_29 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_2_29 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_3_28 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_3_28 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_4_27 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_4_27 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_5_26 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_5_26 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_6_25 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_6_25 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_7_24 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_7_24 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_8_23 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_8_23 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_9_22 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_9_22 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_10_21 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_10_21 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_11_20 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_11_20 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_12_19 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_12_19 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_13_18 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_13_18 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_14_17 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_14_17 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_15_16 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_15_16 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_16_15 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_16_15 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_17_14 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_17_14 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_18_13 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_18_13 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_19_12 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_19_12 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_20_11 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_20_11 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_21_10 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_21_10 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_22_9 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_22_9 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_23_8 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_23_8 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_24_7 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_24_7 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_25_6 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_25_6 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_26_5 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_26_5 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_27_4 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_27_4 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_28_3 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_28_3 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_29_2 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_29_2 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_30_1 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_30_1 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute tilemem_ecp5_inst_0_31_0 MEM_LPC_FILE tilemem_ecp5_inst.lpc
    // exemplar attribute tilemem_ecp5_inst_0_31_0 MEM_INIT_FILE INIT_ALL_0s
    // exemplar end

endmodule
